library verilog;
use verilog.vl_types.all;
entity CLA_testbench is
end CLA_testbench;
