library verilog;
use verilog.vl_types.all;
entity stack_tb is
end stack_tb;
