library verilog;
use verilog.vl_types.all;
entity tb_Lab3_Mealy is
end tb_Lab3_Mealy;
