library verilog;
use verilog.vl_types.all;
entity queue_tb is
end queue_tb;
