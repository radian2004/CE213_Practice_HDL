library verilog;
use verilog.vl_types.all;
entity tb_Lab3_Moore is
end tb_Lab3_Moore;
