library verilog;
use verilog.vl_types.all;
entity locker_tb is
end locker_tb;
